library verilog;
use verilog.vl_types.all;
entity halfAdder_vlg_check_tst is
    port(
        C               : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end halfAdder_vlg_check_tst;
