library verilog;
use verilog.vl_types.all;
entity four_bits_bcd_adder_vlg_check_tst is
    port(
        carry           : in     vl_logic;
        s               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end four_bits_bcd_adder_vlg_check_tst;
