library verilog;
use verilog.vl_types.all;
entity halfAdder_vlg_vec_tst is
end halfAdder_vlg_vec_tst;
