library verilog;
use verilog.vl_types.all;
entity four_bits_bcd_adder_vlg_vec_tst is
end four_bits_bcd_adder_vlg_vec_tst;
