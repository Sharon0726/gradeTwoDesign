library verilog;
use verilog.vl_types.all;
entity fullSub_vlg_vec_tst is
end fullSub_vlg_vec_tst;
