library verilog;
use verilog.vl_types.all;
entity fourBitsBCD_vlg_vec_tst is
end fourBitsBCD_vlg_vec_tst;
