library verilog;
use verilog.vl_types.all;
entity fullSub_vlg_check_tst is
    port(
        Bo              : in     vl_logic;
        Di              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fullSub_vlg_check_tst;
