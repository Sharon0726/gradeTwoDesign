library verilog;
use verilog.vl_types.all;
entity halfSub_vlg_vec_tst is
end halfSub_vlg_vec_tst;
