library verilog;
use verilog.vl_types.all;
entity trippleAdder_vlg_vec_tst is
end trippleAdder_vlg_vec_tst;
